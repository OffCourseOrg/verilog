/*
 *  OffCourse::Verilog
 *		- Home Security UUT
 *
 *  Copyright: Sybe
 *  License: GPLv3 or later
 */

module UUT (

	);


endmodule