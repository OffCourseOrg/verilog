/*
 *  OffCourse::Verilog
 *		- Shift Register DUT
 *
 *  Written by: Sybe
 *  License: MIT
 */

module DUT ();

endmodule