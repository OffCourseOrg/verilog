/*
 *  offcourse::verilog
 *		- ice-cream-mealy UUT
 *
 *  copyright: Aleksandrs
 *  license: GPLv3 or later
 */
 module UUT (
  output wire [?] state
);

endmodule
