/*
 *  OffCourse::Verilog
 *		- Two Wires UUT
 *
 *  Copyright: Sybe
 *  License: GPLv3 or later
 */

module UUT (
		input clk,
		input reset
	);


endmodule