/*
 *  OffCourse::Verilog
 *		- ice-cream-moore UUT
 *
 *  Copyright: Aleksandrs
 *  License: GPLv3 or later
 */

module UUT (

);

endmodule
