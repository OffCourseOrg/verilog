/*
 *  OffCourse::Verilog
 *		- IIC PLACEHOLDER UUT
 *
 *  Copyright: Sybe
 *  License: GPLv3 or later
 */

module UUT (
		input clk,
		input reset
	);


endmodule